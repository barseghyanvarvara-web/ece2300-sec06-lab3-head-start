//========================================================================
// DLatch_GL
//========================================================================

`ifndef DLATCH_GL_V
`define DLATCH_GL_V

// verilator lint_off UNOPTFLAT

module DLatch_GL
(
  input  wire clk,
  input  wire d,
  output wire q
);

  //''' ACTIVITy '''''''''''''''''''''''''''''''''''''''''''''''''''''''''
  // Implement a D Latch using explicit gate-level modeling
  //>'''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

endmodule

// verilator lint_on UNOPTFLAT

`endif /* DLATCH_GL_V */

