//========================================================================
// Register_8b_GL
//========================================================================

`ifndef REGISTER_8B_GL_V
`define REGISTER_8B_GL_V

`include "DFFRE_GL.v"

module Register_8b_GL
(
  input  wire       clk,
  input  wire       rst,
  input  wire       en,
  input  wire [7:0] d,
  output wire [7:0] q
);

  //''' LAB ASSIGNMENT '''''''''''''''''''''''''''''''''''''''''''''''''''
  // Implement an 8-bit register using eight DFFREs
  //>'''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

endmodule

`endif /* REGISTER_8B_GL_V */

