//========================================================================
// DFFRE_GL
//========================================================================

`ifndef DFFRE_GL_V
`define DFFRE_GL_V

`include "DFF_GL.v"
`include "Mux2_1b_GL.v"

// verilator lint_off UNOPTFLAT

module DFFRE_GL
(
  input  wire clk,
  input  wire rst,
  input  wire en,
  input  wire d,
  output wire q
);

  //''' LAB ASSIGNMENT '''''''''''''''''''''''''''''''''''''''''''''''''''
  // Implement a D enabled & resettable flip-flop using DFF and mux
  //>'''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

endmodule

// verilator lint_on UNOPTFLAT

`endif /* DFFRE_GL_V */

