//========================================================================
// Mux2_1b_GL
//========================================================================

`ifndef MUX2_1B_GL
`define MUX2_1B_GL

`include "ece2300/ece2300-misc.v"

module Mux2_1b_GL
(
  (* keep=1 *) input  in0,
  (* keep=1 *) input  in1,
  (* keep=1 *) input  sel,
  (* keep=1 *) output out
);

  //''' LAB ASSIGNMENT '''''''''''''''''''''''''''''''''''''''''''''''''''
  // Implement 1-bit 2-to-1 mux using gate-level modeling
  //>'''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''
  //:
  //: // remove these lines before starting your implementation
  //: `ECE2300_UNUSED( in0 );
  //: `ECE2300_UNUSED( in1 );
  //: `ECE2300_UNUSED( sel );
  //: `ECE2300_UNDRIVEN( out );
  //:

  wire sel_b;
  not( sel_b, sel );

  wire t1;
  and( t1, in0, sel_b );

  wire t2;
  and( t2, in1, sel );

  or( out, t1, t2 );

  //<'''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''

endmodule

`endif /* MUX2_1B_GL */

